module top(a, b, z);
  input a, b;
  output z;
  xor g1 (z, a, b);
endmodule
